// Copyright 2019 © Lockheed Martin Corporation
// Copyright 2019 © Intrinsix Corp.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//    http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
    32'd44, // AIB95ID 63 RX[15]
    32'd45, // AIB95ID 62 RX[14]
    32'd42, // AIB95ID 61 RX[13]
    32'd43, // AIB95ID 60 RX[12]
    32'd40, // AIB95ID 59 RX[11]
    32'd41, // AIB95ID 58 RX[10]
    32'd36, // AIB95ID 57 RX[9]
    32'd37, // AIB95ID 56 RX[8]
    32'd34, // AIB95ID 55 RX[7]
    32'd35, // AIB95ID 54 RX[6]
    32'd32, // AIB95ID 53 RX[5]
    32'd33, // AIB95ID 52 RX[4]
    32'd30, // AIB95ID 51 RX[3]
    32'd31, // AIB95ID 50 RX[2]
    32'd28, // AIB95ID 49 RX[1]
    32'd29, // AIB95ID 48 RX[0]
    32'd27, // AIB95ID 47 SRSTN
    32'd26, // AIB95ID 46 SARSTN
    32'd25, // AIB95ID 45 SPARE[1]
    32'd24, // AIB95ID 44 SPARE[0]
    32'd23, // AIB95ID 43 MARSTN
    32'd22, // AIB95ID 42 MRSTN
    32'd20, // AIB95ID 41 TX[0]
    32'd21, // AIB95ID 40 TX[1]
    32'd18, // AIB95ID 39 TX[2]
    32'd19, // AIB95ID 38 TX[3]
    32'd16, // AIB95ID 37 TX[4]
    32'd17, // AIB95ID 36 TX[5]
    32'd14, // AIB95ID 35 TX[6]
    32'd15, // AIB95ID 34 TX[7]
    32'd12, // AIB95ID 33 TX[8]
    32'd13, // AIB95ID 32 TX[9]
    32'd8 , // AIB95ID 31 TX[10]
    32'd9 , // AIB95ID 30 TX[11]
    32'd6 , // AIB95ID 29 TX[12]
    32'd7 , // AIB95ID 28 TX[13]
    32'd4 , // AIB95ID 27 TX[14]
    32'd5 , // AIB95ID 26 TX[15]
    32'd2 , // AIB95ID 25 TX[16]
    32'd3 , // AIB95ID 24 TX[17]
    32'd0 , // AIB95ID 23 TX[18]
    32'd1 , // AIB95ID 22 TX[19]
    32'd68, // AIB95ID 21 TX[20]
    32'd69, // AIB95ID 20 TX[21]
    32'd66, // AIB95ID 19 TX[22]
    32'd67, // AIB95ID 18 TX[23]
    32'd64, // AIB95ID 17 TX[24]
    32'd65, // AIB95ID 16 TX[25]
    32'd62, // AIB95ID 15 TX[26]
    32'd63, // AIB95ID 14 TX[27]
    32'd60, // AIB95ID 13 TX[28]
    32'd61, // AIB95ID 12 TX[29]
    32'd11, // AIB95ID 11 TXCLKB
    32'd10, // AIB95ID 10 TXCLK
    32'd58, // AIB95ID  9 TX[30]
    32'd59, // AIB95ID  8 TX[31]
    32'd56, // AIB95ID  7 TX[32]
    32'd57, // AIB95ID  6 TX[33]
    32'd54, // AIB95ID  5 TX[34]
    32'd55, // AIB95ID  4 TX[35]
    32'd52, // AIB95ID  3 TX[36]
    32'd53, // AIB95ID  2 TX[37]
    32'd50, // AIB95ID  1 TX[38]
    32'd51  // AIB95ID  0 TX[39]
};
